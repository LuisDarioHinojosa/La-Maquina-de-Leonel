module IntReg(
    input logic [11:0] pc_i,
    input logic c_i,
    input logic z_i,
    input logic clk,
    input logic cen,
    input logic rst,
    input logic we,
    output logic [11:0] pc_o,
    output logic intc_o,
    output logic intz_o
);



logic gateClock;
assign gateClock = clk & cen;	

always_ff @( posedge gateClock ) 
    begin
        if(rst)
            begin
                intc_o <= 0;
                intz_o <= 0;
                pc_o <= 0;
            end
        else if (we)
            begin
                intc_o <= c_i;
                intz_o <= z_i;
                pc_o <= pc_i;
            end
    end

endmodule
