module ALU_GUMNUT(
    input logic [7:0] rs_i,
    input logic [7:0] op2_i,
    input logic [2:0] count_i,
    input logic carry_i,
    input logic [3:0]s_i,
    output logic zero_o,
    output logic carry_o,
    output logic [7:0] res_o

);

endmodule
